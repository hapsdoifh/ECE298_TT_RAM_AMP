magic
tech sky130A
timestamp 1764188770
<< nwell >>
rect 40 160 150 240
rect -100 -20 750 160
<< nmos >>
rect -20 -220 20 -150
rect 170 -220 210 -150
rect 60 -350 130 -310
rect 630 -150 670 -80
rect 480 -290 550 -250
<< pmos >>
rect -20 0 20 140
rect 170 0 210 140
rect 410 0 450 140
rect 630 0 670 140
<< ndiff >>
rect 570 -90 630 -80
rect -80 -160 -20 -150
rect -80 -210 -70 -160
rect -50 -210 -20 -160
rect -80 -220 -20 -210
rect 20 -160 80 -150
rect 20 -210 50 -160
rect 70 -210 80 -160
rect 20 -220 80 -210
rect 110 -160 170 -150
rect 110 -210 120 -160
rect 140 -210 170 -160
rect 110 -220 170 -210
rect 210 -160 270 -150
rect 210 -210 240 -160
rect 260 -210 270 -160
rect 210 -220 270 -210
rect 60 -260 130 -250
rect 60 -280 70 -260
rect 120 -280 130 -260
rect 60 -310 130 -280
rect 60 -380 130 -350
rect 60 -400 70 -380
rect 120 -400 130 -380
rect 60 -410 130 -400
rect 570 -140 580 -90
rect 600 -140 630 -90
rect 570 -150 630 -140
rect 670 -90 730 -80
rect 670 -140 700 -90
rect 720 -140 730 -90
rect 670 -150 730 -140
rect 480 -200 550 -190
rect 480 -220 490 -200
rect 540 -220 550 -200
rect 480 -250 550 -220
rect 480 -320 550 -290
rect 480 -340 490 -320
rect 540 -340 550 -320
rect 480 -350 550 -340
<< pdiff >>
rect -80 130 -20 140
rect -80 10 -70 130
rect -50 10 -20 130
rect -80 0 -20 10
rect 20 130 80 140
rect 20 10 50 130
rect 70 10 80 130
rect 20 0 80 10
rect 110 130 170 140
rect 110 10 120 130
rect 140 10 170 130
rect 110 0 170 10
rect 210 130 270 140
rect 210 10 240 130
rect 260 10 270 130
rect 210 0 270 10
rect 350 130 410 140
rect 350 10 360 130
rect 380 10 410 130
rect 350 0 410 10
rect 450 130 510 140
rect 450 10 480 130
rect 500 10 510 130
rect 450 0 510 10
rect 570 130 630 140
rect 570 10 580 130
rect 600 10 630 130
rect 570 0 630 10
rect 670 130 730 140
rect 670 10 700 130
rect 720 10 730 130
rect 670 0 730 10
<< ndiffc >>
rect -70 -210 -50 -160
rect 50 -210 70 -160
rect 120 -210 140 -160
rect 240 -210 260 -160
rect 70 -280 120 -260
rect 70 -400 120 -380
rect 580 -140 600 -90
rect 700 -140 720 -90
rect 490 -220 540 -200
rect 490 -340 540 -320
<< pdiffc >>
rect -70 10 -50 130
rect 50 10 70 130
rect 120 10 140 130
rect 240 10 260 130
rect 360 10 380 130
rect 480 10 500 130
rect 580 10 600 130
rect 700 10 720 130
<< psubdiff >>
rect 180 -310 260 -290
rect 180 -350 200 -310
rect 240 -350 260 -310
rect 180 -370 260 -350
<< nsubdiff >>
rect 75 205 115 220
rect 75 185 85 205
rect 105 185 115 205
rect 75 170 115 185
<< psubdiffcont >>
rect 200 -350 240 -310
<< nsubdiffcont >>
rect 85 185 105 205
<< poly >>
rect -20 140 20 170
rect 170 140 210 170
rect 410 140 450 170
rect 630 140 670 170
rect -20 -30 20 0
rect -20 -50 -10 -30
rect 10 -50 20 -30
rect -20 -60 20 -50
rect 170 -30 210 0
rect 170 -50 180 -30
rect 200 -50 210 -30
rect 170 -60 210 -50
rect 410 -30 450 0
rect 410 -50 420 -30
rect 440 -50 450 -30
rect 410 -60 450 -50
rect 630 -30 670 0
rect 630 -50 640 -30
rect 660 -50 670 -30
rect 630 -80 670 -50
rect 170 -100 210 -90
rect 170 -120 180 -100
rect 200 -120 210 -100
rect -20 -150 20 -130
rect 170 -150 210 -120
rect -20 -249 20 -220
rect 170 -240 210 -220
rect -20 -269 -11 -249
rect 10 -269 20 -249
rect -20 -280 20 -269
rect 0 -320 60 -310
rect 0 -340 10 -320
rect 30 -340 60 -320
rect 0 -350 60 -340
rect 130 -350 150 -310
rect 630 -170 670 -150
rect 420 -260 480 -250
rect 420 -280 430 -260
rect 450 -280 480 -260
rect 420 -290 480 -280
rect 550 -290 570 -250
<< polycont >>
rect -10 -50 10 -30
rect 180 -50 200 -30
rect 420 -50 440 -30
rect 640 -50 660 -30
rect 180 -120 200 -100
rect -11 -269 10 -249
rect 10 -340 30 -320
rect 430 -280 450 -260
<< xpolycontact >>
rect 330 -410 370 -120
<< locali >>
rect 75 205 115 215
rect 75 185 85 205
rect 105 185 115 205
rect 75 175 115 185
rect -80 130 -40 140
rect -80 10 -70 130
rect -50 10 -40 130
rect -80 0 -40 10
rect 40 130 80 140
rect 40 10 50 130
rect 70 10 80 130
rect 40 0 80 10
rect 110 130 150 140
rect 110 10 120 130
rect 140 10 150 130
rect 110 0 150 10
rect 230 130 270 140
rect 230 10 240 130
rect 260 10 270 130
rect 230 0 270 10
rect 350 130 390 140
rect 350 10 360 130
rect 380 10 390 130
rect -20 -30 20 -20
rect -20 -50 -10 -30
rect 10 -50 20 -30
rect -20 -60 20 -50
rect 170 -30 210 -20
rect 170 -50 180 -30
rect 200 -50 210 -30
rect 170 -60 210 -50
rect 350 -80 390 10
rect 470 130 510 140
rect 470 10 480 130
rect 500 10 510 130
rect 470 0 510 10
rect 570 130 610 140
rect 570 10 580 130
rect 600 10 610 130
rect 570 0 610 10
rect 690 130 730 140
rect 690 10 700 130
rect 720 10 730 130
rect 690 0 730 10
rect 410 -30 450 -20
rect 410 -50 420 -30
rect 440 -50 450 -30
rect 410 -60 450 -50
rect 630 -30 670 -20
rect 630 -50 640 -30
rect 660 -50 670 -30
rect 630 -60 670 -50
rect -140 -100 20 -90
rect -140 -120 -130 -100
rect -110 -120 -10 -100
rect 10 -120 20 -100
rect -140 -130 20 -120
rect 170 -100 210 -90
rect 170 -120 180 -100
rect 200 -120 210 -100
rect 170 -130 210 -120
rect 330 -120 390 -80
rect 570 -90 610 -80
rect 570 -140 580 -90
rect 600 -140 610 -90
rect 570 -150 610 -140
rect 690 -90 730 -80
rect 690 -140 700 -90
rect 720 -140 730 -90
rect 690 -150 730 -140
rect -80 -160 -40 -150
rect -80 -210 -70 -160
rect -50 -210 -40 -160
rect -80 -220 -40 -210
rect 40 -160 80 -150
rect 40 -210 50 -160
rect 70 -210 80 -160
rect 40 -220 80 -210
rect 110 -160 150 -150
rect 110 -210 120 -160
rect 140 -210 150 -160
rect 110 -220 150 -210
rect 230 -160 270 -150
rect 230 -210 240 -160
rect 260 -210 270 -160
rect 230 -220 270 -210
rect -20 -249 20 -240
rect -20 -269 -11 -249
rect 10 -269 20 -249
rect -20 -280 20 -269
rect 60 -260 130 -250
rect 60 -280 70 -260
rect 120 -280 130 -260
rect 60 -290 130 -280
rect 180 -310 260 -290
rect 0 -320 40 -310
rect 0 -340 10 -320
rect 30 -340 40 -320
rect 0 -350 40 -340
rect 180 -350 200 -310
rect 240 -350 260 -310
rect 180 -370 260 -350
rect 480 -200 550 -190
rect 480 -220 490 -200
rect 540 -220 550 -200
rect 480 -230 550 -220
rect 420 -260 460 -250
rect 420 -280 430 -260
rect 450 -280 460 -260
rect 420 -290 460 -280
rect 60 -380 130 -370
rect 60 -400 70 -380
rect 120 -400 130 -380
rect 60 -410 130 -400
rect 480 -320 550 -310
rect 480 -340 490 -320
rect 540 -340 550 -320
rect 480 -350 550 -340
<< viali >>
rect 85 185 105 205
rect -70 10 -50 130
rect 50 10 70 130
rect 120 10 140 130
rect 240 10 260 130
rect 360 10 380 130
rect -10 -50 10 -30
rect 180 -50 200 -30
rect 480 10 500 130
rect 580 10 600 130
rect 700 10 720 130
rect 420 -50 440 -30
rect 640 -50 660 -30
rect -130 -120 -110 -100
rect -10 -120 10 -100
rect 180 -120 200 -100
rect 340 -150 360 -130
rect 580 -140 600 -90
rect 700 -140 720 -90
rect -70 -210 -50 -160
rect 50 -210 70 -160
rect 120 -210 140 -160
rect 240 -210 260 -160
rect -11 -269 10 -249
rect 70 -280 120 -260
rect 10 -340 30 -320
rect 200 -350 240 -310
rect 490 -220 540 -200
rect 430 -280 450 -260
rect 340 -340 360 -320
rect 70 -400 120 -380
rect 490 -340 540 -320
<< metal1 >>
rect -100 240 730 270
rect -140 205 730 240
rect -140 200 85 205
rect 40 185 85 200
rect 105 200 730 205
rect 105 185 150 200
rect 40 160 150 185
rect -80 130 -40 140
rect -80 10 -70 130
rect -50 10 -40 130
rect -80 -20 -40 10
rect 40 130 80 160
rect 40 10 50 130
rect 70 10 80 130
rect 40 0 80 10
rect 110 130 150 160
rect 110 10 120 130
rect 140 10 150 130
rect 110 0 150 10
rect 230 130 270 140
rect 230 10 240 130
rect 260 10 270 130
rect 230 -20 270 10
rect 350 130 390 200
rect 350 10 360 130
rect 380 10 390 130
rect 350 0 390 10
rect 470 130 510 140
rect 470 10 480 130
rect 500 10 510 130
rect -80 -30 210 -20
rect -80 -50 -10 -30
rect 10 -50 180 -30
rect 200 -50 210 -30
rect -80 -60 210 -50
rect 230 -30 450 -20
rect 230 -50 420 -30
rect 440 -50 450 -30
rect 230 -60 450 -50
rect 470 -21 510 10
rect 570 130 610 200
rect 570 10 580 130
rect 600 10 610 130
rect 570 0 610 10
rect 690 130 730 140
rect 690 10 700 130
rect 720 10 730 130
rect 550 -21 670 -20
rect 470 -30 670 -21
rect 470 -50 640 -30
rect 660 -50 670 -30
rect 470 -60 670 -50
rect -140 -100 -100 -90
rect -140 -120 -130 -100
rect -110 -120 -100 -100
rect -140 -130 -100 -120
rect -80 -160 -40 -60
rect -20 -100 210 -90
rect -20 -120 -10 -100
rect 10 -120 180 -100
rect 200 -120 210 -100
rect -20 -130 210 -120
rect -80 -210 -70 -160
rect -50 -210 -40 -160
rect -80 -220 -40 -210
rect 40 -160 80 -150
rect 40 -210 50 -160
rect 70 -180 80 -160
rect 110 -160 150 -150
rect 110 -180 120 -160
rect 70 -210 120 -180
rect 140 -210 150 -160
rect -140 -249 20 -240
rect -140 -269 -11 -249
rect 10 -269 20 -249
rect 40 -250 150 -210
rect 230 -160 270 -60
rect 330 -120 390 -80
rect 330 -130 370 -120
rect 330 -150 340 -130
rect 360 -150 370 -130
rect 330 -160 370 -150
rect 230 -210 240 -160
rect 260 -210 270 -160
rect 230 -220 270 -210
rect 410 -250 450 -60
rect 480 -190 520 -60
rect 570 -90 610 -80
rect 570 -140 580 -90
rect 600 -140 610 -90
rect 480 -200 550 -190
rect 480 -220 490 -200
rect 540 -220 550 -200
rect 480 -230 550 -220
rect -140 -280 20 -269
rect 60 -260 130 -250
rect 60 -280 70 -260
rect 120 -280 130 -260
rect 60 -290 130 -280
rect 410 -260 460 -250
rect 410 -280 430 -260
rect 450 -280 460 -260
rect 410 -290 460 -280
rect 180 -310 260 -290
rect -140 -320 40 -310
rect -140 -340 10 -320
rect 30 -340 40 -320
rect -140 -350 40 -340
rect 180 -350 200 -310
rect 240 -350 260 -310
rect 330 -320 550 -310
rect 330 -340 340 -320
rect 360 -340 490 -320
rect 540 -340 550 -320
rect 330 -350 550 -340
rect 60 -380 130 -370
rect 60 -400 70 -380
rect 120 -400 130 -380
rect 60 -410 130 -400
rect 180 -410 260 -350
rect 570 -410 610 -140
rect 690 -90 730 10
rect 690 -140 700 -90
rect 720 -140 730 -90
rect 690 -150 730 -140
rect -140 -450 610 -410
rect -100 -480 610 -450
<< labels >>
rlabel metal1 55 -40 55 -40 1 VG34
rlabel metal1 -65 235 -64 236 1 Vdd
rlabel viali -120 -110 -120 -110 1 vin2
rlabel metal1 -61 -261 -57 -255 1 vin1
rlabel metal1 90 -450 93 -447 1 Gnd
rlabel metal1 90 -230 90 -230 1 VS12
rlabel metal1 -30 -330 -30 -330 1 Vtail
rlabel metal1 510 -50 520 -40 1 Vout2
rlabel metal1 362 -45 374 -35 1 vinv
rlabel metal1 710 -51 720 -40 1 voutf
rlabel metal1 400 -340 420 -330 1 vbase
<< end >>
